<<<<<<< HEAD
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: D flip flop
// Description: 
// Author: Andy Jeong
//////////////////////////////////////////////////////////////////////////////////

module d_flip_flop(a, b, c);
    output a;
    input b;
    input c;

    reg a;

always @(posedge c)
begin
    a <= b;
end

=======
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: D flip flop
// Description: 
// Author: Andy Jeong
//////////////////////////////////////////////////////////////////////////////////

module d_flip_flop(a, b, c);
    output a;
    input b;
    input c;

    reg a;

always @(posedge c)
begin
    a <= b;
end

>>>>>>> 4c719c418537323adcdba306372967a5ab19167a
endmodule